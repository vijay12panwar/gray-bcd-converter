** GRAY TO BCD CODE CONVERTER**

.subckt inverter 1 2 3
mp 2 1 3 3 pmod w=100u l=1u
mn 2 1 0 0 nmod w=100u l=1u
.model pmod pmos Vt0=-1 kp=80u
.model nmod nmos Vt0=1 kp=200u
.ends

.subckt pass_and 1 2 3 4
m1 1 2 4 4 nmod w=100u l=1u
m2 2 3 4 4 nmod w=100u l=1u
.model nmod nmos Vt0=1 kp=200u
.ends

.subckt pass_or 1 2 3 4
m1 1 3 4 4 nmod w=100u l=1u
m2 2 2 4 4 nmod w=100u l=1u
.model nmod nmos Vt0=1 kp=200u
.ends

Vdd 1 0 dc 5V
Va 10 0 pulse (5 0 0 0 0 32ns 64ns)
Vb 11 0 pulse (5 0 0 0 0 16ns 32ns)
Vc 12 0 pulse (5 0 0 0 0 8ns 16ns)
Vd 13 0 pulse (5 0 0 0 0 4ns 8ns)
xb 10 14 1 inverter
xc 11 15 1 inverter
xd 12 16 1 inverter
xe 13 17 1 inverter
xf 19 35 1 inverter
xg 21 36 1 inverter
xh 22 37 1 inverter
xi 24 38 1 inverter
xj 25 39 1 inverter
xand_one 11 14 10 46 pass_and
xand_two_sub 10 11 15 29 pass_and
xand_two 29 16 12 18 pass_and
xand_three 15 12 16 19 pass_and
x_or_one 18 19 35 47 pass_or
xand_four_suba 14 11 15 30 pass_and
xand_four_subb 30 16 12 31 pass_and
xand_four 31 17 13 20 pass_and
xand_five_suba 15 16 12 32 pass_and
xand_five 32 13 17 21 pass_and
xand_six 10 13 17 22 pass_and
xand_seven_sub 11 12 16 33 pass_and
xor_two_saba 23 21 36 40 pass_or
xor_two_sabb 40 22 37 41 pass_or
xor_two 41 24 38 25 pass_or
xand_seven 33 13 17 23 pass_and
xand_eight_sub 15 12 16 34 pass_and
xand_eight 34 17 13 24 pass_and
xor_three 20 25 39 48 pass_or
.tran 0.1ns 64ns
.control
run
plot V(10)
plot V(11)
plot V(12)
plot V(13)
plot V(10) 
plot V(46) 
plot V(47) 
plot V(48)
.endc
.end